package share_pkg;

integer error_count = 0 ;
integer correct_count = 0 ;
bit test_finsh = 0 ;
    
endpackage

